package SimpleCPU_Parameters;
    typedef int MEM_SIZE;
endpackage:SimpleCPU_Parameters